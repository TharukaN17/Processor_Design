module instr_memory(
    input             clk, write_en,
    input      [15:0] addr, instr_in,
    output reg [15:0] instr_out
    );
    
    reg [15:0] ram [170:0];
    
    parameter loadac    = 8'd4;
    parameter movacr    = 8'd8;
    parameter movacr1   = 8'd9;
    parameter movacr2   = 8'd10;
    parameter movacr3   = 8'd11;
    parameter movacr4   = 8'd12;
    parameter movacr5   = 8'd13;
    parameter movacdar  = 8'd14;
    parameter movrac    = 8'd15;
    parameter movr1ac   = 8'd16;
    parameter movr2ac   = 8'd17;
    parameter movr3ac   = 8'd18;
    parameter movr4ac   = 8'd19;
    parameter movr5ac   = 8'd20;
    parameter movdarac  = 8'd21;
    parameter stac      = 8'd22;
    parameter add       = 8'd25;
    parameter sub       = 8'd27;
    parameter lshift    = 8'd29;
    parameter rshift    = 8'd31;
    parameter incac     = 8'd33;
    parameter incdar    = 8'd34;
    parameter incr1     = 8'd35;
    parameter incr2     = 8'd36;
    parameter incr3     = 8'd37;
    parameter loadim    = 8'd38;
    parameter jumpz     = 8'd41;
    parameter jumpnz    = 8'd48;
    parameter jump      = 8'd49;
    parameter nop       = 8'd50;
    parameter endop     = 8'd51;
    
    initial begin
    ram[0] = loadim;
    ram[1] = 16'd257;
    ram[2] = movacr1;
    ram[3] = movr1ac;
    ram[4] = loadac;
    ram[5] = movacr;
    ram[6] = loadim;
    ram[7] = 8'd2;
    ram[8] = lshift;
    ram[9] = movacr4;
    ram[10] = loadim;
    ram[11] = 8'd1;
    ram[12] = movacr;
    ram[13] = movr1ac;
    ram[14] = add;
    ram[15] = loadac;
    ram[16] = movacr5;
    ram[17] = movr1ac;
    ram[18] = sub;
    ram[19] = loadac;
    ram[20] = movacr;
    ram[21] = movr5ac;
    ram[22] = add;
    ram[23] = movacr5;
    ram[24] = loadim;
    ram[25] = 16'd256;
    ram[26] = movacr;
    ram[27] = movr1ac;
    ram[28] = add;
    ram[29] = loadac;
    ram[30] = movacr;
    ram[31] = movr5ac;
    ram[32] = add;
    ram[33] = movacr5;
    ram[34] = loadim;
    ram[35] = 16'd256;
    ram[36] = movacr;
    ram[37] = movr1ac;
    ram[38] = sub;
    ram[39] = loadac;
    ram[40] = movacr;
    ram[41] = movr5ac;
    ram[42] = add;
    ram[43] = movacr;
    ram[44] = loadim;
    ram[45] = 8'd1;
    ram[46] = lshift;
    ram[47] = movacr;
    ram[48] = movr4ac;
    ram[49] = add;
    ram[50] = movacr4;
    ram[51] = loadim;
    ram[52] = 16'd257;
    ram[53] = movacr;
    ram[54] = movr1ac;
    ram[55] = add;
    ram[56] = loadac;
    ram[57] = movacr5;
    ram[58] = movr1ac;
    ram[59] = sub;
    ram[60] = loadac;
    ram[61] = movacr;
    ram[62] = movr5ac;
    ram[63] = add;
    ram[64] = movacr5;
    ram[65] = loadim;
    ram[66] = 8'd255;
    ram[67] = movacr;
    ram[68] = movr1ac;
    ram[69] = add;
    ram[70] = loadac;
    ram[71] = movacr5;
    ram[72] = movr1ac;
    ram[73] = sub;
    ram[74] = loadac;
    ram[75] = movacr;
    ram[76] = movr5ac;
    ram[77] = add;
    ram[78] = movacr5;
    ram[79] = movacr;
    ram[80] = movr4ac;
    ram[81] = add;
    ram[82] = movacr;
    ram[83] = loadim;
    ram[84] = 8'd4;
    ram[85] = rshift;
    ram[86] = movacr4;
    ram[87] = loadim;
    ram[88] = 16'd257;
    ram[89] = movacr;
    ram[90] = movr1ac;
    ram[91] = sub;
    ram[92] = movacdar;
    ram[93] = movr4ac;
    ram[94] = stac;
    ram[95] = loadim;
    ram[96] = 16'd65278;
    ram[97] = movacr;
    ram[98] = movr1ac;
    ram[99] = sub;
    ram[100] = jumpz;
    ram[101] = 8'd122;
    ram[102] = loadim;
    ram[103] = 8'd253;
    ram[104] = movacr;
    ram[105] = movr2ac;
    ram[106] = sub;
    ram[107] = jumpz;
    ram[108] = 8'd113;
    ram[109] = incr1;
    ram[110] = incr2;
    ram[111] = jump;
    ram[112] = 8'd3;
    ram[113] = incr1;
    ram[114] = incr1;
    ram[115] = incr1;
    ram[116] = loadim;
    ram[117] = 8'd0;
    ram[118] = movacr2;
    ram[119] = jump;
    ram[120] = 8'd3;
    ram[121] = endop;
    ram[122] = loadim;
    ram[123] = 8'd0;
    ram[124] = movacr1; 
    ram[125] = movacr2;
    ram[126] = movacr3;
    ram[127] = movr1ac;
    ram[128] = loadac;
    ram[129] = movacr4;
    ram[130] = movr3ac;
    ram[131] = movacdar; 
    ram[132] = movr4ac;
    ram[133] = stac;
    ram[134] = movr1ac; 
    ram[135] = movacr;
    ram[136] = loadim;
    ram[137] = 16'd64764; 
    ram[138] = sub;
    ram[139] = jumpz;
    ram[140] = 8'd167;
    ram[141] = movr2ac;
    ram[142] = movacr;
    ram[143] = loadim;
    ram[144] = 8'd252;
    ram[145] = sub;
    ram[146] = jumpz;
    ram[147] = 8'd155;
    ram[148] = incr2;
    ram[149] = incr2;
    ram[150] = incr1;
    ram[151] = incr1;
    ram[152] = incr3;
    ram[153] = jump;
    ram[154] = 8'd127;
    ram[155] = loadim;
    ram[156] = 8'd0;
    ram[157] = movacr2;
    ram[158] = loadim;
    ram[159] = 16'd260;
    ram[160] = movacr;
    ram[161] = movr1ac;
    ram[162] = add;
    ram[163] = movacr1;
    ram[164] = incr3;
    ram[165] = jump;
    ram[166] = 8'd127;
    ram[167] = endop;
    end

    always @(posedge clk) begin
        if (write_en == 1)
            ram[addr] <= instr_in;
        else
            instr_out <= ram[addr];
        end
endmodule