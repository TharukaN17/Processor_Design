module instr_memory(
    input             clk, write_en,
    input      [15:0] addr, instr_in,
    output reg [15:0] instr_out
    );
    
    reg [15:0] ram [180:0];
    
    parameter loadac    = 8'd4;
    parameter movacr    = 8'd8;
    parameter movacr1   = 8'd9;
    parameter movacr2   = 8'd10;
    parameter movacr3   = 8'd11;
    parameter movacr4   = 8'd12;
    parameter movacr5   = 8'd13;
    parameter movacdar  = 8'd14;
    parameter movrac    = 8'd15;
    parameter movr1ac   = 8'd16;
    parameter movr2ac   = 8'd17;
    parameter movr3ac   = 8'd18;
    parameter movr4ac   = 8'd19;
    parameter movr5ac   = 8'd20;
    parameter movdarac  = 8'd21;
    parameter stac      = 8'd22;
    parameter add       = 8'd25;
    parameter sub       = 8'd27;
    parameter lshift    = 8'd29;
    parameter rshift    = 8'd31;
    parameter incac     = 8'd33;
    parameter incdar    = 8'd34;
    parameter incr1     = 8'd35;
    parameter incr2     = 8'd36;
    parameter incr3     = 8'd37;
    parameter loadim    = 8'd38;
    parameter jumpz     = 8'd41;
    parameter jumpnz    = 8'd48;
    parameter jump      = 8'd49;
    parameter nop       = 8'd50;
    parameter endop     = 8'd51;
    
    initial begin
    ram[0] = loadim;
    ram[1] = 16'd257;
    ram[2] = movacr1;
    ram[3] = movr1ac;
    ram[4] = loadac;
    ram[5] = movacr;
    ram[6] = loadim;
    ram[7] = 8'd2;
    ram[8] = lshift;
    ram[9] = movacr4;
    ram[10] = loadim;
    ram[11] = 8'd1;
    ram[12] = movacr;
    ram[13] = movr1ac;
    ram[14] = add;
    ram[15] = loadac;
    ram[16] = movacr5;
    ram[17] = movr1ac;
    ram[18] = sub;
    ram[19] = loadac;
    ram[20] = movacr;
    ram[21] = movr5ac;
    ram[22] = add;
    ram[23] = movacr5;
    ram[24] = loadim;
    ram[25] = 16'd256;
    ram[26] = movacr;
    ram[27] = movr1ac;
    ram[28] = add;
    ram[29] = loadac;
    ram[30] = movacr;
    ram[31] = movr5ac;
    ram[32] = add;
    ram[33] = movacr5;
    ram[34] = loadim;
    ram[35] = 16'd256;
    ram[36] = movacr;
    ram[37] = movr1ac;
    ram[38] = sub;
    ram[39] = loadac;
    ram[40] = movacr;
    ram[41] = movr5ac;
    ram[42] = add;
    ram[43] = movacr;
    ram[44] = loadim;
    ram[45] = 8'd1;
    ram[46] = lshift;
    ram[47] = movacr;
    ram[48] = movr4ac;
    ram[49] = add;
    ram[50] = movacr4;
    ram[51] = loadim;
    ram[52] = 16'd257;
    ram[53] = movacr;
    ram[54] = movr1ac;
    ram[55] = add;
    ram[56] = loadac;
    ram[57] = movacr5;
    ram[58] = movr1ac;
    ram[59] = sub;
    ram[60] = loadac;
    ram[61] = movacr;
    ram[62] = movr5ac;
    ram[63] = add;
    ram[64] = movacr5;
    ram[65] = loadim;
    ram[66] = 8'd255;
    ram[67] = movacr;
    ram[68] = movr1ac;
    ram[69] = add;
    ram[70] = loadac;
    ram[71] = movacr;
    ram[72] = movr5ac;
    ram[73] = add;
    ram[74] = movacr5;
    ram[75] = loadim;
    ram[76] = 8'd255;
    ram[77] = movacr;
    ram[78] = movr1ac;
    ram[79] = sub;
    ram[80] = loadac;
    ram[81] = movacr;
    ram[82] = movr5ac;
    ram[83] = add;
    ram[84] = movacr;
    ram[85] = movr4ac;
    ram[86] = add;
    ram[87] = movacr;
    ram[88] = loadim;
    ram[89] = 8'd4;
    ram[90] = rshift;
    ram[91] = movacr4;
    ram[92] = loadim;
    ram[93] = 16'd257;
    ram[94] = movacr;
    ram[95] = movr1ac;
    ram[96] = sub;
    ram[97] = movacdar;
    ram[98] = movr4ac;
    ram[99] = stac;
    ram[100] = loadim;
    ram[101] = 16'd65278;
    ram[102] = movacr;
    ram[103] = movr1ac;
    ram[104] = sub;
    ram[105] = jumpz;
    ram[106] = 8'd127;
    ram[107] = loadim;
    ram[108] = 8'd253;
    ram[109] = movacr;
    ram[110] = movr2ac;
    ram[111] = sub;
    ram[112] = jumpz;
    ram[113] = 8'd118;
    ram[114] = incr1;
    ram[115] = incr2;
    ram[116] = jump;
    ram[117] = 8'd3;
    ram[118] = incr1;
    ram[119] = incr1;
    ram[120] = incr1;
    ram[121] = loadim;
    ram[122] = 8'd0;
    ram[123] = movacr2;
    ram[124] = jump;
    ram[125] = 8'd3;
    ram[126] = endop;
    ram[127] = loadim;
    ram[128] = 8'd0;
    ram[129] = movacr1; 
    ram[130] = movacr2;
    ram[131] = movacr3;
    ram[132] = movr1ac;
    ram[133] = loadac;
    ram[134] = movacr4;
    ram[135] = movr3ac;
    ram[136] = movacdar; 
    ram[137] = movr4ac;
    ram[138] = stac;
    ram[139] = movr1ac; 
    ram[140] = movacr;
    ram[141] = loadim;
    ram[142] = 16'd64764; 
    ram[143] = sub;
    ram[144] = jumpz;
    ram[145] = 8'd172;
    ram[146] = movr2ac;
    ram[147] = movacr;
    ram[148] = loadim;
    ram[149] = 8'd252;
    ram[150] = sub;
    ram[151] = jumpz;
    ram[152] = 8'd160;
    ram[153] = incr2;
    ram[154] = incr2;
    ram[155] = incr1;
    ram[156] = incr1;
    ram[157] = incr3;
    ram[158] = jump;
    ram[159] = 8'd132;
    ram[160] = loadim;
    ram[161] = 8'd0;
    ram[162] = movacr2;
    ram[163] = loadim;
    ram[164] = 16'd260;
    ram[165] = movacr;
    ram[166] = movr1ac;
    ram[167] = add;
    ram[168] = movacr1;
    ram[169] = incr3;
    ram[170] = jump;
    ram[171] = 8'd132;
    ram[172] = endop;
    end

    always @(posedge clk) begin
        if (write_en == 1)
            ram[addr] <= instr_in;
        else
            instr_out <= ram[addr];
        end
endmodule