module instr_memory(
    input             clk, write_en,
    input      [15:0] addr, instr_in,
    output reg [15:0] instr_out
    );
    
    reg [15:0] ram [190:0];
    
    parameter loadac    = 8'd4;
    parameter movacr    = 8'd8;
    parameter movacr1   = 8'd9;
    parameter movacr2   = 8'd10;
    parameter movacr3   = 8'd11;
    parameter movacr4   = 8'd12;
    parameter movacr5   = 8'd13;
    parameter movacdar  = 8'd14;
    parameter movrac    = 8'd15;
    parameter movr1ac   = 8'd16;
    parameter movr2ac   = 8'd17;
    parameter movr3ac   = 8'd18;
    parameter movr4ac   = 8'd19;
    parameter movr5ac   = 8'd20;
    parameter movdarac  = 8'd21;
    parameter stac      = 8'd22;
    parameter add       = 8'd25;
    parameter sub       = 8'd27;
    parameter lshift    = 8'd29;
    parameter rshift    = 8'd31;
    parameter incac     = 8'd33;
    parameter incdar    = 8'd34;
    parameter incr1     = 8'd35;
    parameter incr2     = 8'd36;
    parameter incr3     = 8'd37;
    parameter loadim    = 8'd38;
    parameter jumpz     = 8'd41;
    parameter jumpnz    = 8'd48;
    parameter jump      = 8'd49;
    parameter nop       = 8'd50;
    parameter endop     = 8'd51;
    
    initial begin
    ram[0] = loadim;
    ram[1] = 16'd257; 
    ram[2] = movacr1;
    ram[3] = nop;
    ram[4] = nop; 
    ram[5] = nop;
    ram[6] = nop; 
    ram[7] = nop;
    ram[8] = nop; 
    ram[9] = movr1ac;
    ram[10] = loadac;
    ram[11] = movacr;
    ram[12] = loadim;
    ram[13] = 8'd4;
    ram[14] = lshift;
    ram[15] = movacr4;
    ram[16] = loadim;
    ram[17] = 8'd1;
    ram[18] = movacr;
    ram[19] = movr1ac;
    ram[20] = add;
    ram[21] = loadac;
    ram[22] = movacr5; 
    ram[23] = movr1ac;
    ram[24] = sub ;
    ram[25] = loadac;
    ram[26] = movacr;
    ram[27] = movr5ac;
    ram[28] = add;
    ram[29] = movacr5; 
    ram[30] = loadim;
    ram[31] = 16'd256; 
    ram[32] = movacr;
    ram[33] = movr1ac;
    ram[34] = add;
    ram[35] = loadac;
    ram[36] = movacr;
    ram[37] = movr5ac;
    ram[38] = add;
    ram[39] = movacr5; 
    ram[40] = loadim;
    ram[41] = 16'd256; 
    ram[42] = movacr;
    ram[43] = movr1ac;
    ram[44] = sub;
    ram[45] = loadac;
    ram[46] = movacr;
    ram[47] = movr5ac;
    ram[48] = add;
    ram[49] = movacr5; 
    ram[50] = movacr;
    ram[51] = loadim;
    ram[52] = 8'd1;
    ram[53] = lshift;
    ram[54] = movacr;
    ram[55] = movr5ac;
    ram[56] = add;
    ram[57] = movacr;
    ram[58] = movr4ac;
    ram[59] = add;
    ram[60] = movacr4; 
    ram[61] = loadim;
    ram[62] = 16'd257; 
    ram[63] = movacr;
    ram[64] = movr1ac;
    ram[65] = add;
    ram[66] = loadac;
    ram[67] = movacr5;
    ram[68] = movr1ac;
    ram[69] = sub;
    ram[70] = loadac;
    ram[71] = movacr;
    ram[72] = movr5ac;
    ram[73] = add;
    ram[74] = movacr5;
    ram[75] = loadim;
    ram[76] = 8'd255;
    ram[77] = movacr;
    ram[78] = movr1ac;
    ram[79] = add;
    ram[80] = loadac;
    ram[81] = movacr;
    ram[82] = movr5ac;
    ram[83] = add;
    ram[84] = movacr5;
    ram[85] = loadim;
    ram[86] = 8'd255; 
    ram[87] = movacr;
    ram[88] = movr1ac;
    ram[89] = sub;
    ram[90] = loadac;
    ram[91] = movacr;
    ram[92] = movr5ac;
    ram[93] = add;
    ram[94] = movacr5;
    ram[95] = movacr;
    ram[96] = movr4ac;
    ram[97] = add;
    ram[98] = movacr;
    ram[99] = loadim;
    ram[100] = 8'd5; 
    ram[101] = rshift;
    ram[102] = movacr4;
    ram[103] = loadim;
    ram[104] = 16'd257; 
    ram[105] = movacr;
    ram[106] = movr1ac;
    ram[107] = sub;
    ram[108] = movacdar ;
    ram[109] = movr4ac;
    ram[110] = stac;
    ram[111] = loadim;
    ram[112] = 16'd65278 ; 
    ram[113] = movacr;
    ram[114] = movr1ac;
    ram[115] = sub;
    ram[116] = jumpz;
    ram[117] = 8'd138; 
    ram[118] = loadim;
    ram[119] = 8'd253; 
    ram[120] = movacr;
    ram[121] = movr2ac;
    ram[122] = sub ;
    ram[123] = jumpz;
    ram[124] = 8'd129; 
    ram[125] = incr2; 
    ram[126] = incr1;
    ram[127] = jump;
    ram[128] = 8'd9; 
    ram[129] = incr1;
    ram[130] = incr1;
    ram[131] = incr1;
    ram[132] = loadim;
    ram[133] = 8'd0;
    ram[134] = movacr2;
    ram[135] = jump;
    ram[136] = 8'd9;
    ram[137] = endop; 
    ram[138] = loadim;
    ram[139] = 8'd0;
    ram[140] = movacr1; 
    ram[141] = movacr2;
    ram[142] = movacr3; 
    ram[143] = movr1ac; 
    ram[144] = loadac;
    ram[145] = movacr4;
    ram[146] = movr3ac;
    ram[147] = movacdar ;
    ram[148] = movr4ac;
    ram[149] = stac;
    ram[150] = movr1ac; 
    ram[151] = movacr;
    ram[152] = loadim;
    ram[153] = 16'd64764 ;
    ram[154] = sub;
    ram[155] = jumpz;
    ram[156] = 8'd186;
    ram[157] = movr2ac;
    ram[158] = movacr;
    ram[159] = loadim;
    ram[160] = 8'd252;
    ram[161] = sub;
    ram[162] = jumpz;
    ram[163] = 8'd171;
    ram[164] = incr2;
    ram[165] = incr2;
    ram[166] = incr1;
    ram[167] = incr1;
    ram[168] = incr3;
    ram[169] = jump;
    ram[170] = 8'd143;
    ram[171] = loadim;
    ram[172] = 8'd0;
    ram[173] = movacr2;
    ram[174] = loadim;
    ram[175] = 16'd260;
    ram[176] = movacr;
    ram[177] = movr1ac;
    ram[178] = add;
    ram[179] = movacr1;
    ram[180] = incr3;
    ram[181] = nop;
    ram[182] = nop;
    ram[183] = nop;
    ram[184] = jump;
    ram[185] = 8'd143;
    ram[186] = endop;
    end

    always @(posedge clk) begin
        if (write_en == 1)
            ram[addr] <= instr_in;
        else
            instr_out <= ram[addr];
        end
endmodule